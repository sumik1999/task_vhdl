* /home/kiran99/eSim-Workspace/Subtractor/Subtractor.cir

* EESchema Netlist Version 1.1 (Spice format) creation date: Thu May 13 21:30:58 2021

* To exclude a component from the Spice Netlist add [Spice_Netlist_Enabled] user FIELD set to: N
* To reorder the component spice node sequence add [Spice_Node_Sequence] user FIELD and define sequence: 2,1,0

* Sheet Name: /
U2  A B C Net-_U1-Pad1_ Net-_U1-Pad2_ Net-_U1-Pad3_ adc_bridge_3		
U3  Net-_U1-Pad4_ Net-_U1-Pad5_ DIFF BORROW_OUT dac_bridge_2		
v1  A Net-_R1-Pad2_ pulse		
v2  B Net-_R1-Pad2_ pulse		
v3  C Net-_R1-Pad2_ pulse		
R1  A Net-_R1-Pad2_ 100k		
R2  B Net-_R1-Pad2_ 100k		
R3  C Net-_R1-Pad2_ 100k		
R5  DIFF GND 100k		
R4  BORROW_OUT GND 100k		
U1  Net-_U1-Pad1_ Net-_U1-Pad2_ Net-_U1-Pad3_ Net-_U1-Pad4_ Net-_U1-Pad5_ my_subtractor		

.end
